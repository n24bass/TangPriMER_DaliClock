module data_out
  (
   //
   input wire        clk_lcd,
   output wire [7:0] R,
   output wire [7:0] G,
   output wire [7:0] B,
   input wire        den,
   input wire [10:0] X, // xofs,
   input wire [10:0] Y // yofs
   );

   localparam FONT_START_X = 80; // 188;
   localparam FONT_START_Y = 188;
   localparam FONT_MULTI = 2;
   localparam FONT_HEIGHT = 64 * FONT_MULTI;
   localparam FONT_WIDTH = 45 * FONT_MULTI;
   localparam DOT_WIDTH = 25 * FONT_MULTI;

   reg [7:0]         r_R;
   reg [7:0]         r_G;
   reg [7:0]         r_B;

   reg [5:0]         nframe = 59; // 0..59 60 frame counter

   reg [4:0]         hh;
   reg [4:0]         hh_n;
   reg [5:0]         mm;
   reg [5:0]         mm_n;
   reg [5:0]         ss;
   reg [5:0]         ss_n;

   reg [3:0]         digit; // current digit for dot
   reg [3:0]         digit_n; // next digit 

   reg [5:0]         xofs; // X offset for font
   reg [5:0]         yofs; // Y offset

   reg [5:0]         s[0:3]; // font end poinsts data for digit
   reg [5:0]         f[0:3]; // font end poinsts data for digit_n
   reg [5:0]         ep[0:3]; //

   // functions

   function [23:0] blend_endpoints(
                                   input [5:0] s0, input [5:0] s1, input [5:0] s2, input [5:0] s3, // start
                                   input [5:0] f0, input [5:0] f1, input [5:0] f2, input [5:0] f3, // final
                                   input [7:0] nf // 0..<60 - frame count 
                                   );
      integer                                  i;
      reg [11:0]                               blend;
      reg [11:0]                               v;
      reg [5:0]                                out[0:4];

      // 60 -> 28:32
      localparam MIN = 28;
      localparam MAX = 32;

      begin
         if (nf < MIN) blend = 0;
         else blend = nf - MIN;
         if (MAX < blend) blend = MAX;

         v = ((MAX-blend) * s0 + blend * f0)/MAX;
         out[0] = v[5:0];
         v = ((MAX-blend) * s1 + blend * f1)/MAX;
         out[1] = v[5:0];
         v = ((MAX-blend) * s2 + blend * f2)/MAX;
         out[2] = v[5:0];
         v = ((MAX-blend) * s3 + blend * f3)/MAX;
         out[3] = v[5:0];

         blend_endpoints = {out[0],out[1],out[2],out[3]};
      end
   endfunction // blend_endpoints

   function [24:0] rle_to_endpoints(input [5:0] rle0, input [5:0] rle1, input [5:0] rle2, input [5:0] rle3);
      begin
         if (rle3 != 0)
           rle_to_endpoints = {rle0, rle0 + rle1, rle0 + rle1 + rle2, rle0 + rle1 + rle2 + rle3};
         else
           rle_to_endpoints = {rle0, rle0 + rle1, rle0, rle0 + rle1};
      end
   endfunction // rle_to_endpoints

   function [24:0] font_rle(input [3:0] digit, input [5:0] yofs);
      begin
         case ({digit,yofs})
           // 0
           {4'd0,6'd00}: font_rle = {6'd17,6'd10,6'd00,6'd00};
           {4'd0,6'd01}: font_rle = {6'd15,6'd14,6'd00,6'd00};
           {4'd0,6'd02}: font_rle = {6'd13,6'd07,6'd04,6'd07};
           {4'd0,6'd03}: font_rle = {6'd12,6'd07,6'd06,6'd07};
           {4'd0,6'd04}: font_rle = {6'd11,6'd07,6'd08,6'd07};
           {4'd0,6'd05}: font_rle = {6'd10,6'd07,6'd10,6'd07};
           {4'd0,6'd06}: font_rle = {6'd09,6'd08,6'd10,6'd08};
           {4'd0,6'd07}: font_rle = {6'd08,6'd09,6'd10,6'd09};
           {4'd0,6'd08}: font_rle = {6'd08,6'd08,6'd12,6'd09};
           {4'd0,6'd09}: font_rle = {6'd07,6'd09,6'd12,6'd09};
           {4'd0,6'd10}: font_rle = {6'd06,6'd10,6'd12,6'd10};
           {4'd0,6'd11}: font_rle = {6'd06,6'd10,6'd12,6'd10};
           {4'd0,6'd12}: font_rle = {6'd05,6'd11,6'd12,6'd11};
           {4'd0,6'd13}: font_rle = {6'd05,6'd11,6'd12,6'd11};
           {4'd0,6'd14}: font_rle = {6'd04,6'd12,6'd12,6'd12};
           {4'd0,6'd15}: font_rle = {6'd04,6'd12,6'd12,6'd12};
           {4'd0,6'd16}: font_rle = {6'd04,6'd12,6'd12,6'd12};
           {4'd0,6'd17}: font_rle = {6'd03,6'd13,6'd12,6'd13};
           {4'd0,6'd18}: font_rle = {6'd03,6'd13,6'd13,6'd12};
           {4'd0,6'd19}: font_rle = {6'd03,6'd13,6'd13,6'd12};
           {4'd0,6'd20}: font_rle = {6'd03,6'd13,6'd13,6'd12};
           {4'd0,6'd21}: font_rle = {6'd03,6'd13,6'd13,6'd13};
           {4'd0,6'd22}: font_rle = {6'd02,6'd14,6'd13,6'd13};
           {4'd0,6'd23}: font_rle = {6'd02,6'd14,6'd13,6'd13};
           {4'd0,6'd24}: font_rle = {6'd02,6'd14,6'd13,6'd13};
           {4'd0,6'd25}: font_rle = {6'd02,6'd14,6'd13,6'd13};
           {4'd0,6'd26}: font_rle = {6'd02,6'd14,6'd13,6'd13};
           {4'd0,6'd27}: font_rle = {6'd02,6'd14,6'd13,6'd13};
           {4'd0,6'd28}: font_rle = {6'd02,6'd14,6'd13,6'd13};
           {4'd0,6'd29}: font_rle = {6'd02,6'd14,6'd13,6'd13};
           {4'd0,6'd30}: font_rle = {6'd02,6'd14,6'd13,6'd13};
           {4'd0,6'd31}: font_rle = {6'd02,6'd14,6'd13,6'd13};
           {4'd0,6'd32}: font_rle = {6'd02,6'd14,6'd13,6'd13};
           {4'd0,6'd33}: font_rle = {6'd02,6'd14,6'd13,6'd13};
           {4'd0,6'd34}: font_rle = {6'd02,6'd14,6'd13,6'd13};
           {4'd0,6'd35}: font_rle = {6'd02,6'd14,6'd13,6'd13};
           {4'd0,6'd36}: font_rle = {6'd02,6'd14,6'd13,6'd13};
           {4'd0,6'd37}: font_rle = {6'd02,6'd14,6'd13,6'd13};
           {4'd0,6'd38}: font_rle = {6'd02,6'd14,6'd13,6'd13};
           {4'd0,6'd39}: font_rle = {6'd02,6'd14,6'd13,6'd13};
           {4'd0,6'd40}: font_rle = {6'd02,6'd14,6'd13,6'd13};
           {4'd0,6'd41}: font_rle = {6'd02,6'd14,6'd13,6'd13};
           {4'd0,6'd42}: font_rle = {6'd03,6'd13,6'd13,6'd12};
           {4'd0,6'd43}: font_rle = {6'd03,6'd13,6'd13,6'd12};
           {4'd0,6'd44}: font_rle = {6'd03,6'd13,6'd13,6'd12};
           {4'd0,6'd45}: font_rle = {6'd03,6'd13,6'd12,6'd13};
           {4'd0,6'd46}: font_rle = {6'd04,6'd12,6'd12,6'd12};
           {4'd0,6'd47}: font_rle = {6'd04,6'd12,6'd12,6'd12};
           {4'd0,6'd48}: font_rle = {6'd04,6'd12,6'd12,6'd12};
           {4'd0,6'd49}: font_rle = {6'd05,6'd11,6'd12,6'd11};
           {4'd0,6'd50}: font_rle = {6'd05,6'd11,6'd12,6'd11};
           {4'd0,6'd51}: font_rle = {6'd06,6'd10,6'd12,6'd11};
           {4'd0,6'd52}: font_rle = {6'd06,6'd10,6'd12,6'd10};
           {4'd0,6'd53}: font_rle = {6'd07,6'd09,6'd12,6'd10};
           {4'd0,6'd54}: font_rle = {6'd07,6'd09,6'd12,6'd09};
           {4'd0,6'd55}: font_rle = {6'd08,6'd09,6'd10,6'd09};
           {4'd0,6'd56}: font_rle = {6'd09,6'd08,6'd10,6'd09};
           {4'd0,6'd57}: font_rle = {6'd10,6'd07,6'd10,6'd08};
           {4'd0,6'd58}: font_rle = {6'd10,6'd08,6'd08,6'd08};
           {4'd0,6'd59}: font_rle = {6'd11,6'd07,6'd08,6'd07};
           {4'd0,6'd60}: font_rle = {6'd13,6'd06,6'd06,6'd07};
           {4'd0,6'd61}: font_rle = {6'd14,6'd07,6'd02,6'd07};
           {4'd0,6'd62}: font_rle = {6'd16,6'd12,6'd00,6'd00};
           {4'd0,6'd63}: font_rle = {6'd19,6'd06,6'd00,6'd00};
           // 1
           {4'd1,6'd00}: font_rle = {6'd26,6'd04,6'd00,6'd00};
           {4'd1,6'd01}: font_rle = {6'd24,6'd06,6'd00,6'd00};
           {4'd1,6'd02}: font_rle = {6'd22,6'd08,6'd00,6'd00};
           {4'd1,6'd03}: font_rle = {6'd19,6'd11,6'd00,6'd00};
           {4'd1,6'd04}: font_rle = {6'd17,6'd13,6'd00,6'd00};
           {4'd1,6'd05}: font_rle = {6'd15,6'd15,6'd00,6'd00};
           {4'd1,6'd06}: font_rle = {6'd12,6'd18,6'd00,6'd00};
           {4'd1,6'd07}: font_rle = {6'd10,6'd20,6'd00,6'd00};
           {4'd1,6'd08}: font_rle = {6'd08,6'd22,6'd00,6'd00};
           {4'd1,6'd09}: font_rle = {6'd05,6'd25,6'd00,6'd00};
           {4'd1,6'd10}: font_rle = {6'd05,6'd03,6'd07,6'd15};
           {4'd1,6'd11}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd12}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd13}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd14}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd15}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd16}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd17}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd18}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd19}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd20}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd21}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd22}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd23}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd24}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd25}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd26}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd27}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd28}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd29}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd30}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd31}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd32}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd33}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd34}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd35}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd36}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd37}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd38}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd39}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd40}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd41}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd42}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd43}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd44}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd45}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd46}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd47}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd48}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd49}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd50}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd51}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd52}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd53}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd54}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd55}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd56}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd57}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd1,6'd58}: font_rle = {6'd15,6'd16,6'd00,6'd00};
           {4'd1,6'd59}: font_rle = {6'd15,6'd16,6'd00,6'd00};
           {4'd1,6'd60}: font_rle = {6'd13,6'd19,6'd00,6'd00};
           {4'd1,6'd61}: font_rle = {6'd11,6'd23,6'd00,6'd00};
           {4'd1,6'd62}: font_rle = {6'd05,6'd35,6'd00,6'd00};
           {4'd1,6'd63}: font_rle = {6'd05,6'd35,6'd00,6'd00};
           // 2
           {4'd2,6'd00}: font_rle = {6'd17,6'd12,6'd00,6'd00};
           {4'd2,6'd01}: font_rle = {6'd15,6'd16,6'd00,6'd00};
           {4'd2,6'd02}: font_rle = {6'd13,6'd20,6'd00,6'd00};
           {4'd2,6'd03}: font_rle = {6'd12,6'd22,6'd00,6'd00};
           {4'd2,6'd04}: font_rle = {6'd11,6'd24,6'd00,6'd00};
           {4'd2,6'd05}: font_rle = {6'd09,6'd27,6'd00,6'd00};
           {4'd2,6'd06}: font_rle = {6'd09,6'd28,6'd00,6'd00};
           {4'd2,6'd07}: font_rle = {6'd08,6'd30,6'd00,6'd00};
           {4'd2,6'd08}: font_rle = {6'd07,6'd31,6'd00,6'd00};
           {4'd2,6'd09}: font_rle = {6'd06,6'd33,6'd00,6'd00};
           {4'd2,6'd10}: font_rle = {6'd06,6'd06,6'd08,6'd19};
           {4'd2,6'd11}: font_rle = {6'd05,6'd05,6'd12,6'd17};
           {4'd2,6'd12}: font_rle = {6'd05,6'd04,6'd15,6'd16};
           {4'd2,6'd13}: font_rle = {6'd04,6'd04,6'd17,6'd15};
           {4'd2,6'd14}: font_rle = {6'd04,6'd03,6'd18,6'd15};
           {4'd2,6'd15}: font_rle = {6'd03,6'd03,6'd20,6'd14};
           {4'd2,6'd16}: font_rle = {6'd03,6'd03,6'd20,6'd14};
           {4'd2,6'd17}: font_rle = {6'd03,6'd02,6'd22,6'd13};
           {4'd2,6'd18}: font_rle = {6'd27,6'd13,6'd00,6'd00};
           {4'd2,6'd19}: font_rle = {6'd27,6'd13,6'd00,6'd00};
           {4'd2,6'd20}: font_rle = {6'd27,6'd13,6'd00,6'd00};
           {4'd2,6'd21}: font_rle = {6'd27,6'd13,6'd00,6'd00};
           {4'd2,6'd22}: font_rle = {6'd28,6'd11,6'd00,6'd00};
           {4'd2,6'd23}: font_rle = {6'd27,6'd12,6'd00,6'd00};
           {4'd2,6'd24}: font_rle = {6'd27,6'd12,6'd00,6'd00};
           {4'd2,6'd25}: font_rle = {6'd27,6'd11,6'd00,6'd00};
           {4'd2,6'd26}: font_rle = {6'd27,6'd11,6'd00,6'd00};
           {4'd2,6'd27}: font_rle = {6'd27,6'd10,6'd00,6'd00};
           {4'd2,6'd28}: font_rle = {6'd26,6'd10,6'd00,6'd00};
           {4'd2,6'd29}: font_rle = {6'd26,6'd10,6'd00,6'd00};
           {4'd2,6'd30}: font_rle = {6'd26,6'd09,6'd00,6'd00};
           {4'd2,6'd31}: font_rle = {6'd25,6'd09,6'd00,6'd00};
           {4'd2,6'd32}: font_rle = {6'd25,6'd09,6'd00,6'd00};
           {4'd2,6'd33}: font_rle = {6'd24,6'd09,6'd00,6'd00};
           {4'd2,6'd34}: font_rle = {6'd24,6'd08,6'd00,6'd00};
           {4'd2,6'd35}: font_rle = {6'd23,6'd08,6'd00,6'd00};
           {4'd2,6'd36}: font_rle = {6'd22,6'd08,6'd00,6'd00};
           {4'd2,6'd37}: font_rle = {6'd22,6'd07,6'd00,6'd00};
           {4'd2,6'd38}: font_rle = {6'd21,6'd07,6'd00,6'd00};
           {4'd2,6'd39}: font_rle = {6'd20,6'd07,6'd00,6'd00};
           {4'd2,6'd40}: font_rle = {6'd20,6'd06,6'd00,6'd00};
           {4'd2,6'd41}: font_rle = {6'd19,6'd06,6'd00,6'd00};
           {4'd2,6'd42}: font_rle = {6'd18,6'd06,6'd00,6'd00};
           {4'd2,6'd43}: font_rle = {6'd17,6'd05,6'd00,6'd00};
           {4'd2,6'd44}: font_rle = {6'd16,6'd05,6'd00,6'd00};
           {4'd2,6'd45}: font_rle = {6'd16,6'd04,6'd21,6'd03};
           {4'd2,6'd46}: font_rle = {6'd15,6'd04,6'd22,6'd02};
           {4'd2,6'd47}: font_rle = {6'd14,6'd04,6'd22,6'd03};
           {4'd2,6'd48}: font_rle = {6'd13,6'd04,6'd23,6'd03};
           {4'd2,6'd49}: font_rle = {6'd12,6'd04,6'd23,6'd04};
           {4'd2,6'd50}: font_rle = {6'd11,6'd04,6'd23,6'd04};
           {4'd2,6'd51}: font_rle = {6'd10,6'd05,6'd19,6'd08};
           {4'd2,6'd52}: font_rle = {6'd10,6'd32,6'd00,6'd00};
           {4'd2,6'd53}: font_rle = {6'd09,6'd33,6'd00,6'd00};
           {4'd2,6'd54}: font_rle = {6'd08,6'd34,6'd00,6'd00};
           {4'd2,6'd55}: font_rle = {6'd07,6'd34,6'd00,6'd00};
           {4'd2,6'd56}: font_rle = {6'd06,6'd35,6'd00,6'd00};
           {4'd2,6'd57}: font_rle = {6'd05,6'd36,6'd00,6'd00};
           {4'd2,6'd58}: font_rle = {6'd04,6'd37,6'd00,6'd00};
           {4'd2,6'd59}: font_rle = {6'd03,6'd38,6'd00,6'd00};
           {4'd2,6'd60}: font_rle = {6'd02,6'd38,6'd00,6'd00};
           {4'd2,6'd61}: font_rle = {6'd01,6'd39,6'd00,6'd00};
           {4'd2,6'd62}: font_rle = {6'd01,6'd39,6'd00,6'd00};
           {4'd2,6'd63}: font_rle = {6'd01,6'd39,6'd00,6'd00};   
           // 3
           {4'd3,6'd00}: font_rle = {6'd18,6'd12,6'd00,6'd00};
           {4'd3,6'd01}: font_rle = {6'd15,6'd17,6'd00,6'd00};
           {4'd3,6'd02}: font_rle = {6'd13,6'd21,6'd00,6'd00};
           {4'd3,6'd03}: font_rle = {6'd12,6'd23,6'd00,6'd00};
           {4'd3,6'd04}: font_rle = {6'd10,6'd26,6'd00,6'd00};
           {4'd3,6'd05}: font_rle = {6'd09,6'd28,6'd00,6'd00};
           {4'd3,6'd06}: font_rle = {6'd08,6'd30,6'd00,6'd00};
           {4'd3,6'd07}: font_rle = {6'd07,6'd05,6'd09,6'd17};
           {4'd3,6'd08}: font_rle = {6'd06,6'd04,6'd12,6'd16};
           {4'd3,6'd09}: font_rle = {6'd06,6'd03,6'd15,6'd15};
           {4'd3,6'd10}: font_rle = {6'd05,6'd03,6'd16,6'd15};
           {4'd3,6'd11}: font_rle = {6'd04,6'd03,6'd18,6'd14};
           {4'd3,6'd12}: font_rle = {6'd04,6'd02,6'd19,6'd14};
           {4'd3,6'd13}: font_rle = {6'd04,6'd02,6'd20,6'd13};
           {4'd3,6'd14}: font_rle = {6'd26,6'd13,6'd00,6'd00};
           {4'd3,6'd15}: font_rle = {6'd26,6'd13,6'd00,6'd00};
           {4'd3,6'd16}: font_rle = {6'd26,6'd12,6'd00,6'd00};
           {4'd3,6'd17}: font_rle = {6'd26,6'd12,6'd00,6'd00};
           {4'd3,6'd18}: font_rle = {6'd26,6'd11,6'd00,6'd00};
           {4'd3,6'd19}: font_rle = {6'd26,6'd11,6'd00,6'd00};
           {4'd3,6'd20}: font_rle = {6'd25,6'd11,6'd00,6'd00};
           {4'd3,6'd21}: font_rle = {6'd25,6'd10,6'd00,6'd00};
           {4'd3,6'd22}: font_rle = {6'd24,6'd09,6'd00,6'd00};
           {4'd3,6'd23}: font_rle = {6'd23,6'd09,6'd00,6'd00};
           {4'd3,6'd24}: font_rle = {6'd22,6'd11,6'd00,6'd00};
           {4'd3,6'd25}: font_rle = {6'd21,6'd14,6'd00,6'd00};
           {4'd3,6'd26}: font_rle = {6'd19,6'd17,6'd00,6'd00};
           {4'd3,6'd27}: font_rle = {6'd17,6'd21,6'd00,6'd00};
           {4'd3,6'd28}: font_rle = {6'd14,6'd25,6'd00,6'd00};
           {4'd3,6'd29}: font_rle = {6'd14,6'd25,6'd00,6'd00};
           {4'd3,6'd30}: font_rle = {6'd16,6'd24,6'd00,6'd00};
           {4'd3,6'd31}: font_rle = {6'd19,6'd22,6'd00,6'd00};
           {4'd3,6'd32}: font_rle = {6'd21,6'd20,6'd00,6'd00};
           {4'd3,6'd33}: font_rle = {6'd23,6'd18,6'd00,6'd00};
           {4'd3,6'd34}: font_rle = {6'd24,6'd18,6'd00,6'd00};
           {4'd3,6'd35}: font_rle = {6'd26,6'd16,6'd00,6'd00};
           {4'd3,6'd36}: font_rle = {6'd27,6'd15,6'd00,6'd00};
           {4'd3,6'd37}: font_rle = {6'd28,6'd14,6'd00,6'd00};
           {4'd3,6'd38}: font_rle = {6'd29,6'd14,6'd00,6'd00};
           {4'd3,6'd39}: font_rle = {6'd30,6'd13,6'd00,6'd00};
           {4'd3,6'd40}: font_rle = {6'd30,6'd13,6'd00,6'd00};
           {4'd3,6'd41}: font_rle = {6'd31,6'd12,6'd00,6'd00};
           {4'd3,6'd42}: font_rle = {6'd31,6'd11,6'd00,6'd00};
           {4'd3,6'd43}: font_rle = {6'd32,6'd10,6'd00,6'd00};
           {4'd3,6'd44}: font_rle = {6'd32,6'd10,6'd00,6'd00};
           {4'd3,6'd45}: font_rle = {6'd32,6'd10,6'd00,6'd00};
           {4'd3,6'd46}: font_rle = {6'd32,6'd10,6'd00,6'd00};
           {4'd3,6'd47}: font_rle = {6'd33,6'd08,6'd00,6'd00};
           {4'd3,6'd48}: font_rle = {6'd33,6'd08,6'd00,6'd00};
           {4'd3,6'd49}: font_rle = {6'd33,6'd08,6'd00,6'd00};
           {4'd3,6'd50}: font_rle = {6'd05,6'd04,6'd23,6'd08};
           {4'd3,6'd51}: font_rle = {6'd03,6'd08,6'd21,6'd07};
           {4'd3,6'd52}: font_rle = {6'd02,6'd11,6'd19,6'd07};
           {4'd3,6'd53}: font_rle = {6'd02,6'd12,6'd18,6'd06};
           {4'd3,6'd54}: font_rle = {6'd01,6'd14,6'd16,6'd06};
           {4'd3,6'd55}: font_rle = {6'd01,6'd15,6'd15,6'd05};
           {4'd3,6'd56}: font_rle = {6'd01,6'd16,6'd13,6'd05};
           {4'd3,6'd57}: font_rle = {6'd02,6'd16,6'd11,6'd05};
           {4'd3,6'd58}: font_rle = {6'd02,6'd18,6'd08,6'd05};
           {4'd3,6'd59}: font_rle = {6'd03,6'd19,6'd03,6'd06};
           {4'd3,6'd60}: font_rle = {6'd03,6'd27,6'd00,6'd00};
           {4'd3,6'd61}: font_rle = {6'd05,6'd23,6'd00,6'd00};
           {4'd3,6'd62}: font_rle = {6'd07,6'd18,6'd00,6'd00};
           {4'd3,6'd63}: font_rle = {6'd11,6'd09,6'd00,6'd00};
           // 4
           {4'd4,6'd00}: font_rle = {6'd30,6'd08,6'd00,6'd00};
           {4'd4,6'd01}: font_rle = {6'd29,6'd09,6'd00,6'd00};
           {4'd4,6'd02}: font_rle = {6'd28,6'd10,6'd00,6'd00};
           {4'd4,6'd03}: font_rle = {6'd27,6'd11,6'd00,6'd00};
           {4'd4,6'd04}: font_rle = {6'd27,6'd11,6'd00,6'd00};
           {4'd4,6'd05}: font_rle = {6'd26,6'd12,6'd00,6'd00};
           {4'd4,6'd06}: font_rle = {6'd25,6'd13,6'd00,6'd00};
           {4'd4,6'd07}: font_rle = {6'd24,6'd14,6'd00,6'd00};
           {4'd4,6'd08}: font_rle = {6'd24,6'd14,6'd00,6'd00};
           {4'd4,6'd09}: font_rle = {6'd23,6'd15,6'd00,6'd00};
           {4'd4,6'd10}: font_rle = {6'd22,6'd16,6'd00,6'd00};
           {4'd4,6'd11}: font_rle = {6'd21,6'd17,6'd00,6'd00};
           {4'd4,6'd12}: font_rle = {6'd20,6'd18,6'd00,6'd00};
           {4'd4,6'd13}: font_rle = {6'd20,6'd18,6'd00,6'd00};
           {4'd4,6'd14}: font_rle = {6'd19,6'd19,6'd00,6'd00};
           {4'd4,6'd15}: font_rle = {6'd18,6'd05,6'd01,6'd14};
           {4'd4,6'd16}: font_rle = {6'd17,6'd05,6'd02,6'd14};
           {4'd4,6'd17}: font_rle = {6'd17,6'd04,6'd03,6'd14};
           {4'd4,6'd18}: font_rle = {6'd16,6'd04,6'd04,6'd14};
           {4'd4,6'd19}: font_rle = {6'd15,6'd05,6'd04,6'd14};
           {4'd4,6'd20}: font_rle = {6'd14,6'd05,6'd05,6'd14};
           {4'd4,6'd21}: font_rle = {6'd14,6'd04,6'd06,6'd14};
           {4'd4,6'd22}: font_rle = {6'd13,6'd05,6'd06,6'd14};
           {4'd4,6'd23}: font_rle = {6'd12,6'd05,6'd07,6'd14};
           {4'd4,6'd24}: font_rle = {6'd12,6'd04,6'd08,6'd14};
           {4'd4,6'd25}: font_rle = {6'd11,6'd04,6'd09,6'd14};
           {4'd4,6'd26}: font_rle = {6'd10,6'd05,6'd09,6'd14};
           {4'd4,6'd27}: font_rle = {6'd09,6'd05,6'd10,6'd14};
           {4'd4,6'd28}: font_rle = {6'd09,6'd04,6'd11,6'd14};
           {4'd4,6'd29}: font_rle = {6'd08,6'd04,6'd12,6'd14};
           {4'd4,6'd30}: font_rle = {6'd07,6'd05,6'd12,6'd14};
           {4'd4,6'd31}: font_rle = {6'd07,6'd04,6'd13,6'd14};
           {4'd4,6'd32}: font_rle = {6'd06,6'd04,6'd14,6'd14};
           {4'd4,6'd33}: font_rle = {6'd05,6'd05,6'd14,6'd14};
           {4'd4,6'd34}: font_rle = {6'd05,6'd04,6'd15,6'd14};
           {4'd4,6'd35}: font_rle = {6'd04,6'd04,6'd16,6'd14};
           {4'd4,6'd36}: font_rle = {6'd03,6'd04,6'd17,6'd14};
           {4'd4,6'd37}: font_rle = {6'd02,6'd05,6'd17,6'd14};
           {4'd4,6'd38}: font_rle = {6'd02,6'd04,6'd18,6'd14};
           {4'd4,6'd39}: font_rle = {6'd01,6'd04,6'd19,6'd14};
           {4'd4,6'd40}: font_rle = {6'd01,6'd42,6'd00,6'd00};
           {4'd4,6'd41}: font_rle = {6'd01,6'd42,6'd00,6'd00};
           {4'd4,6'd42}: font_rle = {6'd01,6'd42,6'd00,6'd00};
           {4'd4,6'd43}: font_rle = {6'd01,6'd42,6'd00,6'd00};
           {4'd4,6'd44}: font_rle = {6'd01,6'd42,6'd00,6'd00};
           {4'd4,6'd45}: font_rle = {6'd01,6'd42,6'd00,6'd00};
           {4'd4,6'd46}: font_rle = {6'd01,6'd42,6'd00,6'd00};
           {4'd4,6'd47}: font_rle = {6'd01,6'd42,6'd00,6'd00};
           {4'd4,6'd48}: font_rle = {6'd01,6'd42,6'd00,6'd00};
           {4'd4,6'd49}: font_rle = {6'd01,6'd42,6'd00,6'd00};
           {4'd4,6'd50}: font_rle = {6'd24,6'd14,6'd00,6'd00};
           {4'd4,6'd51}: font_rle = {6'd24,6'd14,6'd00,6'd00};
           {4'd4,6'd52}: font_rle = {6'd24,6'd14,6'd00,6'd00};
           {4'd4,6'd53}: font_rle = {6'd24,6'd14,6'd00,6'd00};
           {4'd4,6'd54}: font_rle = {6'd24,6'd14,6'd00,6'd00};
           {4'd4,6'd55}: font_rle = {6'd24,6'd14,6'd00,6'd00};
           {4'd4,6'd56}: font_rle = {6'd24,6'd14,6'd00,6'd00};
           {4'd4,6'd57}: font_rle = {6'd24,6'd14,6'd00,6'd00};
           {4'd4,6'd58}: font_rle = {6'd24,6'd14,6'd00,6'd00};
           {4'd4,6'd59}: font_rle = {6'd24,6'd14,6'd00,6'd00};
           {4'd4,6'd60}: font_rle = {6'd24,6'd14,6'd00,6'd00};
           {4'd4,6'd61}: font_rle = {6'd24,6'd14,6'd00,6'd00};
           {4'd4,6'd62}: font_rle = {6'd24,6'd14,6'd00,6'd00};
           {4'd4,6'd63}: font_rle = {6'd24,6'd14,6'd00,6'd00};
           // 5
           {4'd5,6'd00}: font_rle = {6'd13,6'd30,6'd00,6'd00};
           {4'd5,6'd01}: font_rle = {6'd13,6'd30,6'd00,6'd00};
           {4'd5,6'd02}: font_rle = {6'd13,6'd30,6'd00,6'd00};
           {4'd5,6'd03}: font_rle = {6'd13,6'd29,6'd00,6'd00};
           {4'd5,6'd04}: font_rle = {6'd12,6'd30,6'd00,6'd00};
           {4'd5,6'd05}: font_rle = {6'd12,6'd30,6'd00,6'd00};
           {4'd5,6'd06}: font_rle = {6'd12,6'd29,6'd00,6'd00};
           {4'd5,6'd07}: font_rle = {6'd11,6'd30,6'd00,6'd00};
           {4'd5,6'd08}: font_rle = {6'd11,6'd30,6'd00,6'd00};
           {4'd5,6'd09}: font_rle = {6'd11,6'd29,6'd00,6'd00};
           {4'd5,6'd10}: font_rle = {6'd11,6'd29,6'd00,6'd00};
           {4'd5,6'd11}: font_rle = {6'd10,6'd04,6'd00,6'd00};
           {4'd5,6'd12}: font_rle = {6'd10,6'd03,6'd00,6'd00};
           {4'd5,6'd13}: font_rle = {6'd10,6'd03,6'd00,6'd00};
           {4'd5,6'd14}: font_rle = {6'd10,6'd03,6'd00,6'd00};
           {4'd5,6'd15}: font_rle = {6'd09,6'd03,6'd00,6'd00};
           {4'd5,6'd16}: font_rle = {6'd09,6'd03,6'd00,6'd00};
           {4'd5,6'd17}: font_rle = {6'd09,6'd03,6'd00,6'd00};
           {4'd5,6'd18}: font_rle = {6'd08,6'd04,6'd00,6'd00};
           {4'd5,6'd19}: font_rle = {6'd08,6'd07,6'd00,6'd00};
           {4'd5,6'd20}: font_rle = {6'd08,6'd15,6'd00,6'd00};
           {4'd5,6'd21}: font_rle = {6'd08,6'd19,6'd00,6'd00};
           {4'd5,6'd22}: font_rle = {6'd07,6'd22,6'd00,6'd00};
           {4'd5,6'd23}: font_rle = {6'd07,6'd25,6'd00,6'd00};
           {4'd5,6'd24}: font_rle = {6'd07,6'd26,6'd00,6'd00};
           {4'd5,6'd25}: font_rle = {6'd06,6'd29,6'd00,6'd00};
           {4'd5,6'd26}: font_rle = {6'd06,6'd30,6'd00,6'd00};
           {4'd5,6'd27}: font_rle = {6'd06,6'd31,6'd00,6'd00};
           {4'd5,6'd28}: font_rle = {6'd06,6'd32,6'd00,6'd00};
           {4'd5,6'd29}: font_rle = {6'd05,6'd34,6'd00,6'd00};
           {4'd5,6'd30}: font_rle = {6'd05,6'd34,6'd00,6'd00};
           {4'd5,6'd31}: font_rle = {6'd05,6'd35,6'd00,6'd00};
           {4'd5,6'd32}: font_rle = {6'd13,6'd27,6'd00,6'd00};
           {4'd5,6'd33}: font_rle = {6'd19,6'd22,6'd00,6'd00};
           {4'd5,6'd34}: font_rle = {6'd22,6'd19,6'd00,6'd00};
           {4'd5,6'd35}: font_rle = {6'd24,6'd17,6'd00,6'd00};
           {4'd5,6'd36}: font_rle = {6'd26,6'd16,6'd00,6'd00};
           {4'd5,6'd37}: font_rle = {6'd28,6'd14,6'd00,6'd00};
           {4'd5,6'd38}: font_rle = {6'd29,6'd13,6'd00,6'd00};
           {4'd5,6'd39}: font_rle = {6'd31,6'd11,6'd00,6'd00};
           {4'd5,6'd40}: font_rle = {6'd32,6'd10,6'd00,6'd00};
           {4'd5,6'd41}: font_rle = {6'd33,6'd09,6'd00,6'd00};
           {4'd5,6'd42}: font_rle = {6'd33,6'd09,6'd00,6'd00};
           {4'd5,6'd43}: font_rle = {6'd34,6'd08,6'd00,6'd00};
           {4'd5,6'd44}: font_rle = {6'd34,6'd08,6'd00,6'd00};
           {4'd5,6'd45}: font_rle = {6'd35,6'd07,6'd00,6'd00};
           {4'd5,6'd46}: font_rle = {6'd35,6'd06,6'd00,6'd00};
           {4'd5,6'd47}: font_rle = {6'd35,6'd06,6'd00,6'd00};
           {4'd5,6'd48}: font_rle = {6'd35,6'd06,6'd00,6'd00};
           {4'd5,6'd49}: font_rle = {6'd35,6'd05,6'd00,6'd00};
           {4'd5,6'd50}: font_rle = {6'd05,6'd05,6'd25,6'd05};
           {4'd5,6'd51}: font_rle = {6'd04,6'd08,6'd23,6'd04};
           {4'd5,6'd52}: font_rle = {6'd03,6'd11,6'd20,6'd05};
           {4'd5,6'd53}: font_rle = {6'd02,6'd14,6'd18,6'd04};
           {4'd5,6'd54}: font_rle = {6'd02,6'd15,6'd16,6'd04};
           {4'd5,6'd55}: font_rle = {6'd02,6'd16,6'd14,6'd05};
           {4'd5,6'd56}: font_rle = {6'd02,6'd18,6'd11,6'd05};
           {4'd5,6'd57}: font_rle = {6'd02,6'd20,6'd08,6'd04};
           {4'd5,6'd58}: font_rle = {6'd03,6'd30,6'd00,6'd00};
           {4'd5,6'd59}: font_rle = {6'd03,6'd29,6'd00,6'd00};
           {4'd5,6'd60}: font_rle = {6'd04,6'd26,6'd00,6'd00};
           {4'd5,6'd61}: font_rle = {6'd06,6'd22,6'd00,6'd00};
           {4'd5,6'd62}: font_rle = {6'd08,6'd17,6'd00,6'd00};
           {4'd5,6'd63}: font_rle = {6'd11,6'd09,6'd00,6'd00};
           // 6
           {4'd6,6'd00}: font_rle = {6'd36,6'd07,6'd00,6'd00};
           {4'd6,6'd01}: font_rle = {6'd32,6'd10,6'd00,6'd00};
           {4'd6,6'd02}: font_rle = {6'd29,6'd10,6'd00,6'd00};
           {4'd6,6'd03}: font_rle = {6'd26,6'd10,6'd00,6'd00};
           {4'd6,6'd04}: font_rle = {6'd24,6'd10,6'd00,6'd00};
           {4'd6,6'd05}: font_rle = {6'd22,6'd10,6'd00,6'd00};
           {4'd6,6'd06}: font_rle = {6'd20,6'd10,6'd00,6'd00};
           {4'd6,6'd07}: font_rle = {6'd19,6'd10,6'd00,6'd00};
           {4'd6,6'd08}: font_rle = {6'd17,6'd11,6'd00,6'd00};
           {4'd6,6'd09}: font_rle = {6'd16,6'd11,6'd00,6'd00};
           {4'd6,6'd10}: font_rle = {6'd15,6'd11,6'd00,6'd00};
           {4'd6,6'd11}: font_rle = {6'd13,6'd12,6'd00,6'd00};
           {4'd6,6'd12}: font_rle = {6'd12,6'd12,6'd00,6'd00};
           {4'd6,6'd13}: font_rle = {6'd11,6'd12,6'd00,6'd00};
           {4'd6,6'd14}: font_rle = {6'd11,6'd11,6'd00,6'd00};
           {4'd6,6'd15}: font_rle = {6'd10,6'd12,6'd00,6'd00};
           {4'd6,6'd16}: font_rle = {6'd09,6'd12,6'd00,6'd00};
           {4'd6,6'd17}: font_rle = {6'd08,6'd13,6'd00,6'd00};
           {4'd6,6'd18}: font_rle = {6'd08,6'd12,6'd00,6'd00};
           {4'd6,6'd19}: font_rle = {6'd07,6'd13,6'd00,6'd00};
           {4'd6,6'd20}: font_rle = {6'd06,6'd13,6'd00,6'd00};
           {4'd6,6'd21}: font_rle = {6'd06,6'd13,6'd00,6'd00};
           {4'd6,6'd22}: font_rle = {6'd05,6'd14,6'd00,6'd00};
           {4'd6,6'd23}: font_rle = {6'd05,6'd13,6'd00,6'd00};
           {4'd6,6'd24}: font_rle = {6'd05,6'd13,6'd04,6'd08};
           {4'd6,6'd25}: font_rle = {6'd04,6'd29,6'd00,6'd00};
           {4'd6,6'd26}: font_rle = {6'd04,6'd31,6'd00,6'd00};
           {4'd6,6'd27}: font_rle = {6'd04,6'd33,6'd00,6'd00};
           {4'd6,6'd28}: font_rle = {6'd03,6'd15,6'd06,6'd14};
           {4'd6,6'd29}: font_rle = {6'd03,6'd14,6'd09,6'd13};
           {4'd6,6'd30}: font_rle = {6'd03,6'd14,6'd09,6'd14};
           {4'd6,6'd31}: font_rle = {6'd03,6'd14,6'd10,6'd13};
           {4'd6,6'd32}: font_rle = {6'd03,6'd14,6'd11,6'd13};
           {4'd6,6'd33}: font_rle = {6'd02,6'd14,6'd12,6'd13};
           {4'd6,6'd34}: font_rle = {6'd02,6'd14,6'd12,6'd14};
           {4'd6,6'd35}: font_rle = {6'd02,6'd14,6'd12,6'd14};
           {4'd6,6'd36}: font_rle = {6'd02,6'd14,6'd13,6'd13};
           {4'd6,6'd37}: font_rle = {6'd02,6'd14,6'd13,6'd14};
           {4'd6,6'd38}: font_rle = {6'd02,6'd14,6'd13,6'd14};
           {4'd6,6'd39}: font_rle = {6'd02,6'd14,6'd13,6'd14};
           {4'd6,6'd40}: font_rle = {6'd02,6'd14,6'd13,6'd14};
           {4'd6,6'd41}: font_rle = {6'd02,6'd14,6'd13,6'd14};
           {4'd6,6'd42}: font_rle = {6'd02,6'd14,6'd13,6'd14};
           {4'd6,6'd43}: font_rle = {6'd03,6'd13,6'd13,6'd14};
           {4'd6,6'd44}: font_rle = {6'd03,6'd13,6'd13,6'd14};
           {4'd6,6'd45}: font_rle = {6'd03,6'd13,6'd13,6'd14};
           {4'd6,6'd46}: font_rle = {6'd03,6'd13,6'd13,6'd14};
           {4'd6,6'd47}: font_rle = {6'd03,6'd13,6'd13,6'd14};
           {4'd6,6'd48}: font_rle = {6'd04,6'd12,6'd13,6'd13};
           {4'd6,6'd49}: font_rle = {6'd04,6'd13,6'd12,6'd13};
           {4'd6,6'd50}: font_rle = {6'd04,6'd13,6'd12,6'd13};
           {4'd6,6'd51}: font_rle = {6'd05,6'd12,6'd12,6'd12};
           {4'd6,6'd52}: font_rle = {6'd05,6'd12,6'd12,6'd12};
           {4'd6,6'd53}: font_rle = {6'd06,6'd11,6'd12,6'd12};
           {4'd6,6'd54}: font_rle = {6'd06,6'd11,6'd12,6'd11};
           {4'd6,6'd55}: font_rle = {6'd07,6'd10,6'd12,6'd10};
           {4'd6,6'd56}: font_rle = {6'd08,6'd10,6'd11,6'd10};
           {4'd6,6'd57}: font_rle = {6'd09,6'd09,6'd11,6'd09};
           {4'd6,6'd58}: font_rle = {6'd10,6'd09,6'd09,6'd09};
           {4'd6,6'd59}: font_rle = {6'd11,6'd08,6'd09,6'd08};
           {4'd6,6'd60}: font_rle = {6'd12,6'd08,6'd07,6'd07};
           {4'd6,6'd61}: font_rle = {6'd14,6'd08,6'd03,6'd08};
           {4'd6,6'd62}: font_rle = {6'd16,6'd14,6'd00,6'd00};
           {4'd6,6'd63}: font_rle = {6'd19,6'd08,6'd00,6'd00};
           // 7
           {4'd7,6'd00}: font_rle = {6'd05,6'd39,6'd00,6'd00};
           {4'd7,6'd01}: font_rle = {6'd04,6'd39,6'd00,6'd00};
           {4'd7,6'd02}: font_rle = {6'd04,6'd39,6'd00,6'd00};
           {4'd7,6'd03}: font_rle = {6'd04,6'd39,6'd00,6'd00};
           {4'd7,6'd04}: font_rle = {6'd04,6'd38,6'd00,6'd00};
           {4'd7,6'd05}: font_rle = {6'd04,6'd38,6'd00,6'd00};
           {4'd7,6'd06}: font_rle = {6'd03,6'd39,6'd00,6'd00};
           {4'd7,6'd07}: font_rle = {6'd03,6'd38,6'd00,6'd00};
           {4'd7,6'd08}: font_rle = {6'd03,6'd38,6'd00,6'd00};
           {4'd7,6'd09}: font_rle = {6'd03,6'd38,6'd00,6'd00};
           {4'd7,6'd10}: font_rle = {6'd03,6'd37,6'd00,6'd00};
           {4'd7,6'd11}: font_rle = {6'd02,6'd38,6'd00,6'd00};
           {4'd7,6'd12}: font_rle = {6'd02,6'd08,6'd21,6'd08};
           {4'd7,6'd13}: font_rle = {6'd02,6'd05,6'd24,6'd08};
           {4'd7,6'd14}: font_rle = {6'd02,6'd03,6'd26,6'd08};
           {4'd7,6'd15}: font_rle = {6'd02,6'd03,6'd26,6'd07};
           {4'd7,6'd16}: font_rle = {6'd01,6'd03,6'd26,6'd08};
           {4'd7,6'd17}: font_rle = {6'd01,6'd03,6'd26,6'd08};
           {4'd7,6'd18}: font_rle = {6'd01,6'd02,6'd27,6'd07};
           {4'd7,6'd19}: font_rle = {6'd01,6'd02,6'd26,6'd08};
           {4'd7,6'd20}: font_rle = {6'd29,6'd08,6'd00,6'd00};
           {4'd7,6'd21}: font_rle = {6'd29,6'd07,6'd00,6'd00};
           {4'd7,6'd22}: font_rle = {6'd28,6'd08,6'd00,6'd00};
           {4'd7,6'd23}: font_rle = {6'd28,6'd08,6'd00,6'd00};
           {4'd7,6'd24}: font_rle = {6'd27,6'd08,6'd00,6'd00};
           {4'd7,6'd25}: font_rle = {6'd27,6'd08,6'd00,6'd00};
           {4'd7,6'd26}: font_rle = {6'd27,6'd08,6'd00,6'd00};
           {4'd7,6'd27}: font_rle = {6'd26,6'd08,6'd00,6'd00};
           {4'd7,6'd28}: font_rle = {6'd26,6'd08,6'd00,6'd00};
           {4'd7,6'd29}: font_rle = {6'd26,6'd08,6'd00,6'd00};
           {4'd7,6'd30}: font_rle = {6'd25,6'd08,6'd00,6'd00};
           {4'd7,6'd31}: font_rle = {6'd25,6'd08,6'd00,6'd00};
           {4'd7,6'd32}: font_rle = {6'd25,6'd08,6'd00,6'd00};
           {4'd7,6'd33}: font_rle = {6'd24,6'd08,6'd00,6'd00};
           {4'd7,6'd34}: font_rle = {6'd24,6'd08,6'd00,6'd00};
           {4'd7,6'd35}: font_rle = {6'd23,6'd08,6'd00,6'd00};
           {4'd7,6'd36}: font_rle = {6'd23,6'd08,6'd00,6'd00};
           {4'd7,6'd37}: font_rle = {6'd23,6'd08,6'd00,6'd00};
           {4'd7,6'd38}: font_rle = {6'd22,6'd08,6'd00,6'd00};
           {4'd7,6'd39}: font_rle = {6'd22,6'd08,6'd00,6'd00};
           {4'd7,6'd40}: font_rle = {6'd22,6'd08,6'd00,6'd00};
           {4'd7,6'd41}: font_rle = {6'd21,6'd08,6'd00,6'd00};
           {4'd7,6'd42}: font_rle = {6'd21,6'd08,6'd00,6'd00};
           {4'd7,6'd43}: font_rle = {6'd20,6'd09,6'd00,6'd00};
           {4'd7,6'd44}: font_rle = {6'd20,6'd08,6'd00,6'd00};
           {4'd7,6'd45}: font_rle = {6'd20,6'd08,6'd00,6'd00};
           {4'd7,6'd46}: font_rle = {6'd19,6'd09,6'd00,6'd00};
           {4'd7,6'd47}: font_rle = {6'd19,6'd08,6'd00,6'd00};
           {4'd7,6'd48}: font_rle = {6'd19,6'd08,6'd00,6'd00};
           {4'd7,6'd49}: font_rle = {6'd18,6'd09,6'd00,6'd00};
           {4'd7,6'd50}: font_rle = {6'd18,6'd08,6'd00,6'd00};
           {4'd7,6'd51}: font_rle = {6'd18,6'd08,6'd00,6'd00};
           {4'd7,6'd52}: font_rle = {6'd17,6'd09,6'd00,6'd00};
           {4'd7,6'd53}: font_rle = {6'd17,6'd08,6'd00,6'd00};
           {4'd7,6'd54}: font_rle = {6'd16,6'd09,6'd00,6'd00};
           {4'd7,6'd55}: font_rle = {6'd16,6'd09,6'd00,6'd00};
           {4'd7,6'd56}: font_rle = {6'd16,6'd08,6'd00,6'd00};
           {4'd7,6'd57}: font_rle = {6'd15,6'd09,6'd00,6'd00};
           {4'd7,6'd58}: font_rle = {6'd15,6'd09,6'd00,6'd00};
           {4'd7,6'd59}: font_rle = {6'd15,6'd08,6'd00,6'd00};
           {4'd7,6'd60}: font_rle = {6'd14,6'd09,6'd00,6'd00};
           {4'd7,6'd61}: font_rle = {6'd14,6'd08,6'd00,6'd00};
           {4'd7,6'd62}: font_rle = {6'd14,6'd08,6'd00,6'd00};
           {4'd7,6'd63}: font_rle = {6'd13,6'd09,6'd00,6'd00};
           // 8
           {4'd8,6'd00}: font_rle = {6'd16,6'd15,6'd00,6'd00};
           {4'd8,6'd01}: font_rle = {6'd13,6'd21,6'd00,6'd00};
           {4'd8,6'd02}: font_rle = {6'd11,6'd08,6'd07,6'd10};
           {4'd8,6'd03}: font_rle = {6'd10,6'd07,6'd10,6'd10};
           {4'd8,6'd04}: font_rle = {6'd08,6'd08,6'd12,6'd10};
           {4'd8,6'd05}: font_rle = {6'd07,6'd09,6'd13,6'd10};
           {4'd8,6'd06}: font_rle = {6'd06,6'd09,6'd14,6'd11};
           {4'd8,6'd07}: font_rle = {6'd05,6'd10,6'd15,6'd10};
           {4'd8,6'd08}: font_rle = {6'd05,6'd10,6'd15,6'd11};
           {4'd8,6'd09}: font_rle = {6'd04,6'd11,6'd15,6'd11};
           {4'd8,6'd10}: font_rle = {6'd04,6'd11,6'd15,6'd11};
           {4'd8,6'd11}: font_rle = {6'd04,6'd11,6'd16,6'd10};
           {4'd8,6'd12}: font_rle = {6'd03,6'd12,6'd16,6'd10};
           {4'd8,6'd13}: font_rle = {6'd03,6'd12,6'd16,6'd10};
           {4'd8,6'd14}: font_rle = {6'd03,6'd13,6'd15,6'd10};
           {4'd8,6'd15}: font_rle = {6'd03,6'd13,6'd15,6'd10};
           {4'd8,6'd16}: font_rle = {6'd03,6'd14,6'd13,6'd11};
           {4'd8,6'd17}: font_rle = {6'd03,6'd15,6'd12,6'd10};
           {4'd8,6'd18}: font_rle = {6'd03,6'd16,6'd11,6'd09};
           {4'd8,6'd19}: font_rle = {6'd03,6'd17,6'd10,6'd09};
           {4'd8,6'd20}: font_rle = {6'd04,6'd17,6'd08,6'd09};
           {4'd8,6'd21}: font_rle = {6'd04,6'd18,6'd06,6'd09};
           {4'd8,6'd22}: font_rle = {6'd05,6'd19,6'd04,6'd07};
           {4'd8,6'd23}: font_rle = {6'd05,6'd21,6'd01,6'd06};
           {4'd8,6'd24}: font_rle = {6'd06,6'd25,6'd00,6'd00};
           {4'd8,6'd25}: font_rle = {6'd07,6'd22,6'd00,6'd00};
           {4'd8,6'd26}: font_rle = {6'd07,6'd23,6'd00,6'd00};
           {4'd8,6'd27}: font_rle = {6'd08,6'd23,6'd00,6'd00};
           {4'd8,6'd28}: font_rle = {6'd10,6'd23,6'd00,6'd00};
           {4'd8,6'd29}: font_rle = {6'd11,6'd23,6'd00,6'd00};
           {4'd8,6'd30}: font_rle = {6'd12,6'd23,6'd00,6'd00};
           {4'd8,6'd31}: font_rle = {6'd13,6'd23,6'd00,6'd00};
           {4'd8,6'd32}: font_rle = {6'd15,6'd22,6'd00,6'd00};
           {4'd8,6'd33}: font_rle = {6'd15,6'd23,6'd00,6'd00};
           {4'd8,6'd34}: font_rle = {6'd12,6'd27,6'd00,6'd00};
           {4'd8,6'd35}: font_rle = {6'd10,6'd07,6'd02,6'd21};
           {4'd8,6'd36}: font_rle = {6'd08,6'd08,6'd05,6'd19};
           {4'd8,6'd37}: font_rle = {6'd07,6'd09,6'd06,6'd19};
           {4'd8,6'd38}: font_rle = {6'd06,6'd09,6'd08,6'd18};
           {4'd8,6'd39}: font_rle = {6'd05,6'd09,6'd11,6'd17};
           {4'd8,6'd40}: font_rle = {6'd04,6'd10,6'd12,6'd16};
           {4'd8,6'd41}: font_rle = {6'd04,6'd10,6'd13,6'd15};
           {4'd8,6'd42}: font_rle = {6'd03,6'd10,6'd14,6'd15};
           {4'd8,6'd43}: font_rle = {6'd03,6'd10,6'd15,6'd14};
           {4'd8,6'd44}: font_rle = {6'd02,6'd11,6'd16,6'd13};
           {4'd8,6'd45}: font_rle = {6'd02,6'd11,6'd16,6'd13};
           {4'd8,6'd46}: font_rle = {6'd02,6'd11,6'd16,6'd13};
           {4'd8,6'd47}: font_rle = {6'd02,6'd11,6'd17,6'd12};
           {4'd8,6'd48}: font_rle = {6'd02,6'd11,6'd17,6'd12};
           {4'd8,6'd49}: font_rle = {6'd02,6'd11,6'd17,6'd12};
           {4'd8,6'd50}: font_rle = {6'd02,6'd11,6'd17,6'd12};
           {4'd8,6'd51}: font_rle = {6'd02,6'd11,6'd17,6'd12};
           {4'd8,6'd52}: font_rle = {6'd03,6'd10,6'd17,6'd11};
           {4'd8,6'd53}: font_rle = {6'd03,6'd10,6'd17,6'd11};
           {4'd8,6'd54}: font_rle = {6'd03,6'd11,6'd16,6'd10};
           {4'd8,6'd55}: font_rle = {6'd04,6'd10,6'd15,6'd11};
           {4'd8,6'd56}: font_rle = {6'd04,6'd10,6'd15,6'd10};
           {4'd8,6'd57}: font_rle = {6'd05,6'd10,6'd14,6'd09};
           {4'd8,6'd58}: font_rle = {6'd06,6'd10,6'd12,6'd09};
           {4'd8,6'd59}: font_rle = {6'd07,6'd10,6'd10,6'd09};
           {4'd8,6'd60}: font_rle = {6'd09,6'd09,6'd07,6'd09};
           {4'd8,6'd61}: font_rle = {6'd11,6'd21,6'd00,6'd00};
           {4'd8,6'd62}: font_rle = {6'd13,6'd17,6'd00,6'd00};
           {4'd8,6'd63}: font_rle = {6'd17,6'd09,6'd00,6'd00};
           // 9
           {4'd9,6'd00}: font_rle = {6'd16,6'd12,6'd00,6'd00};
           {4'd9,6'd01}: font_rle = {6'd13,6'd17,6'd00,6'd00};
           {4'd9,6'd02}: font_rle = {6'd11,6'd08,6'd05,6'd08};
           {4'd9,6'd03}: font_rle = {6'd10,6'd08,6'd07,6'd09};
           {4'd9,6'd04}: font_rle = {6'd09,6'd08,6'd09,6'd09};
           {4'd9,6'd05}: font_rle = {6'd08,6'd09,6'd10,6'd09};
           {4'd9,6'd06}: font_rle = {6'd07,6'd09,6'd11,6'd10};
           {4'd9,6'd07}: font_rle = {6'd06,6'd10,6'd11,6'd10};
           {4'd9,6'd08}: font_rle = {6'd05,6'd11,6'd12,6'd10};
           {4'd9,6'd09}: font_rle = {6'd05,6'd11,6'd12,6'd11};
           {4'd9,6'd10}: font_rle = {6'd04,6'd11,6'd13,6'd11};
           {4'd9,6'd11}: font_rle = {6'd04,6'd11,6'd13,6'd12};
           {4'd9,6'd12}: font_rle = {6'd03,6'd12,6'd13,6'd12};
           {4'd9,6'd13}: font_rle = {6'd03,6'd12,6'd13,6'd13};
           {4'd9,6'd14}: font_rle = {6'd03,6'd12,6'd14,6'd12};
           {4'd9,6'd15}: font_rle = {6'd03,6'd12,6'd14,6'd12};
           {4'd9,6'd16}: font_rle = {6'd02,6'd13,6'd14,6'd13};
           {4'd9,6'd17}: font_rle = {6'd02,6'd13,6'd14,6'd13};
           {4'd9,6'd18}: font_rle = {6'd02,6'd13,6'd14,6'd13};
           {4'd9,6'd19}: font_rle = {6'd02,6'd13,6'd14,6'd13};
           {4'd9,6'd20}: font_rle = {6'd02,6'd13,6'd14,6'd13};
           {4'd9,6'd21}: font_rle = {6'd02,6'd14,6'd13,6'd14};
           {4'd9,6'd22}: font_rle = {6'd02,6'd14,6'd13,6'd14};
           {4'd9,6'd23}: font_rle = {6'd02,6'd14,6'd13,6'd14};
           {4'd9,6'd24}: font_rle = {6'd02,6'd14,6'd13,6'd14};
           {4'd9,6'd25}: font_rle = {6'd03,6'd13,6'd13,6'd14};
           {4'd9,6'd26}: font_rle = {6'd03,6'd13,6'd13,6'd14};
           {4'd9,6'd27}: font_rle = {6'd03,6'd13,6'd13,6'd14};
           {4'd9,6'd28}: font_rle = {6'd03,6'd14,6'd12,6'd14};
           {4'd9,6'd29}: font_rle = {6'd04,6'd13,6'd12,6'd14};
           {4'd9,6'd30}: font_rle = {6'd04,6'd13,6'd12,6'd13};
           {4'd9,6'd31}: font_rle = {6'd05,6'd13,6'd10,6'd14};
           {4'd9,6'd32}: font_rle = {6'd05,6'd13,6'd10,6'd14};
           {4'd9,6'd33}: font_rle = {6'd06,6'd13,6'd09,6'd14};
           {4'd9,6'd34}: font_rle = {6'd07,6'd13,6'd08,6'd14};
           {4'd9,6'd35}: font_rle = {6'd08,6'd15,6'd01,6'd17};
           {4'd9,6'd36}: font_rle = {6'd09,6'd32,6'd00,6'd00};
           {4'd9,6'd37}: font_rle = {6'd11,6'd30,6'd00,6'd00};
           {4'd9,6'd38}: font_rle = {6'd13,6'd11,6'd03,6'd14};
           {4'd9,6'd39}: font_rle = {6'd27,6'd13,6'd00,6'd00};
           {4'd9,6'd40}: font_rle = {6'd26,6'd14,6'd00,6'd00};
           {4'd9,6'd41}: font_rle = {6'd26,6'd13,6'd00,6'd00};
           {4'd9,6'd42}: font_rle = {6'd26,6'd13,6'd00,6'd00};
           {4'd9,6'd43}: font_rle = {6'd25,6'd13,6'd00,6'd00};
           {4'd9,6'd44}: font_rle = {6'd25,6'd13,6'd00,6'd00};
           {4'd9,6'd45}: font_rle = {6'd25,6'd12,6'd00,6'd00};
           {4'd9,6'd46}: font_rle = {6'd24,6'd12,6'd00,6'd00};
           {4'd9,6'd47}: font_rle = {6'd24,6'd12,6'd00,6'd00};
           {4'd9,6'd48}: font_rle = {6'd23,6'd12,6'd00,6'd00};
           {4'd9,6'd49}: font_rle = {6'd22,6'd12,6'd00,6'd00};
           {4'd9,6'd50}: font_rle = {6'd22,6'd11,6'd00,6'd00};
           {4'd9,6'd51}: font_rle = {6'd21,6'd11,6'd00,6'd00};
           {4'd9,6'd52}: font_rle = {6'd20,6'd11,6'd00,6'd00};
           {4'd9,6'd53}: font_rle = {6'd19,6'd11,6'd00,6'd00};
           {4'd9,6'd54}: font_rle = {6'd18,6'd10,6'd00,6'd00};
           {4'd9,6'd55}: font_rle = {6'd17,6'd10,6'd00,6'd00};
           {4'd9,6'd56}: font_rle = {6'd16,6'd10,6'd00,6'd00};
           {4'd9,6'd57}: font_rle = {6'd14,6'd10,6'd00,6'd00};
           {4'd9,6'd58}: font_rle = {6'd12,6'd10,6'd00,6'd00};
           {4'd9,6'd59}: font_rle = {6'd10,6'd10,6'd00,6'd00};
           {4'd9,6'd60}: font_rle = {6'd08,6'd10,6'd00,6'd00};
           {4'd9,6'd61}: font_rle = {6'd04,6'd11,6'd00,6'd00};
           {4'd9,6'd62}: font_rle = {6'd03,6'd08,6'd00,6'd00};
           {4'd9,6'd63}: font_rle = {6'd03,6'd03,6'd00,6'd00};
           // :
           {4'd10,6'd00}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd10,6'd01}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd10,6'd02}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd10,6'd03}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd10,6'd04}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd10,6'd05}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd10,6'd06}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd10,6'd07}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd10,6'd08}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd10,6'd09}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd10,6'd10}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd10,6'd11}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd10,6'd12}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd10,6'd13}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd10,6'd14}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd10,6'd15}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd10,6'd16}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd10,6'd17}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd10,6'd18}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd10,6'd19}: font_rle = {6'd09,6'd07,6'd00,6'd00};
           {4'd10,6'd20}: font_rle = {6'd08,6'd10,6'd00,6'd00};
           {4'd10,6'd21}: font_rle = {6'd07,6'd12,6'd00,6'd00};
           {4'd10,6'd22}: font_rle = {6'd06,6'd13,6'd00,6'd00};
           {4'd10,6'd23}: font_rle = {6'd06,6'd14,6'd00,6'd00};
           {4'd10,6'd24}: font_rle = {6'd06,6'd14,6'd00,6'd00};
           {4'd10,6'd25}: font_rle = {6'd05,6'd15,6'd00,6'd00};
           {4'd10,6'd26}: font_rle = {6'd05,6'd15,6'd00,6'd00};
           {4'd10,6'd27}: font_rle = {6'd05,6'd15,6'd00,6'd00};
           {4'd10,6'd28}: font_rle = {6'd06,6'd14,6'd00,6'd00};
           {4'd10,6'd29}: font_rle = {6'd06,6'd14,6'd00,6'd00};
           {4'd10,6'd30}: font_rle = {6'd06,6'd13,6'd00,6'd00};
           {4'd10,6'd31}: font_rle = {6'd07,6'd12,6'd00,6'd00};
           {4'd10,6'd32}: font_rle = {6'd08,6'd10,6'd00,6'd00};
           {4'd10,6'd33}: font_rle = {6'd10,6'd06,6'd00,6'd00};
           {4'd10,6'd34}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd10,6'd35}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd10,6'd36}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd10,6'd37}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd10,6'd38}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd10,6'd39}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd10,6'd40}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd10,6'd41}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd10,6'd42}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd10,6'd43}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd10,6'd44}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd10,6'd45}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd10,6'd46}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd10,6'd47}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd10,6'd48}: font_rle = {6'd12,6'd02,6'd00,6'd00};
           {4'd10,6'd49}: font_rle = {6'd09,6'd08,6'd00,6'd00};
           {4'd10,6'd50}: font_rle = {6'd08,6'd10,6'd00,6'd00};
           {4'd10,6'd51}: font_rle = {6'd07,6'd12,6'd00,6'd00};
           {4'd10,6'd52}: font_rle = {6'd06,6'd14,6'd00,6'd00};
           {4'd10,6'd53}: font_rle = {6'd06,6'd14,6'd00,6'd00};
           {4'd10,6'd54}: font_rle = {6'd05,6'd15,6'd00,6'd00};
           {4'd10,6'd55}: font_rle = {6'd05,6'd15,6'd00,6'd00};
           {4'd10,6'd56}: font_rle = {6'd05,6'd15,6'd00,6'd00};
           {4'd10,6'd57}: font_rle = {6'd05,6'd15,6'd00,6'd00};
           {4'd10,6'd58}: font_rle = {6'd06,6'd14,6'd00,6'd00};
           {4'd10,6'd59}: font_rle = {6'd06,6'd14,6'd00,6'd00};
           {4'd10,6'd60}: font_rle = {6'd07,6'd12,6'd00,6'd00};
           {4'd10,6'd61}: font_rle = {6'd07,6'd11,6'd00,6'd00};
           {4'd10,6'd62}: font_rle = {6'd09,6'd08,6'd00,6'd00};
           {4'd10,6'd63}: font_rle = {6'd11,6'd04,6'd00,6'd00};
           // -
           {4'd11,6'd00}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd01}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd02}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd03}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd04}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd05}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd06}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd07}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd08}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd09}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd10}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd11}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd12}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd13}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd14}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd15}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd16}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd17}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd18}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd19}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd20}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd21}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd22}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd23}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd24}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd25}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd26}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd27}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd28}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd29}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd30}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd31}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd32}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd33}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd34}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd35}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd36}: font_rle = {6'd02,6'd21,6'd00,6'd00};
           {4'd11,6'd37}: font_rle = {6'd02,6'd21,6'd00,6'd00};
           {4'd11,6'd38}: font_rle = {6'd02,6'd21,6'd00,6'd00};
           {4'd11,6'd39}: font_rle = {6'd02,6'd21,6'd00,6'd00};
           {4'd11,6'd40}: font_rle = {6'd02,6'd21,6'd00,6'd00};
           {4'd11,6'd41}: font_rle = {6'd02,6'd21,6'd00,6'd00};
           {4'd11,6'd42}: font_rle = {6'd02,6'd21,6'd00,6'd00};
           {4'd11,6'd43}: font_rle = {6'd02,6'd21,6'd00,6'd00};
           {4'd11,6'd44}: font_rle = {6'd02,6'd21,6'd00,6'd00};
           {4'd11,6'd45}: font_rle = {6'd02,6'd21,6'd00,6'd00};
           {4'd11,6'd46}: font_rle = {6'd02,6'd21,6'd00,6'd00};
           {4'd11,6'd47}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd48}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd49}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd50}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd51}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd52}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd53}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd54}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd55}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd56}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd57}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd58}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd59}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd60}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd61}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd62}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           {4'd11,6'd63}: font_rle = {6'd32,6'd00,6'd00,6'd00};
           //
           default: font_rle = {6'd00,6'd00,6'd00,6'd00};
         endcase // case (caseexpr)
      end
   endfunction

   function [16:0] incr_hms(input [4:0] h, input [5:0] m, input [5:0] s);
      begin
         s = s + 1;
         if (60 <= s) begin
            s = 0;
            m = m + 1;
            if (60 <= m) begin
               m = 0;
               h = h + 1;
               if (24 <= h) begin
                  h = 0;
               end
            end
         end
         
         incr_hms = {h,m,s};
      end
   endfunction // incr_hms

   // --

   initial begin
      {hh,mm,ss} = {5'd15, 6'd10, 6'd0}; // initial value
      {hh_n,mm_n,ss_n} = incr_hms(hh,mm,ss);
   end
   
   // --

   // `define BLINK_COLON
   
   always@(posedge clk_lcd) begin
      if (den) begin
         if (X == 0 && Y == 0) nframe = nframe + 1;
         if (nframe >= 60) begin
            nframe = 0;
            {hh,mm,ss} = {hh_n,mm_n,ss_n};
            {hh_n,mm_n,ss_n} = incr_hms(hh,mm,ss);
         end

         if (FONT_START_Y <= Y && Y < FONT_START_Y + FONT_HEIGHT) begin
            yofs = (Y - FONT_START_Y) / FONT_MULTI;

            if (FONT_START_X <= X && X < FONT_START_X + FONT_WIDTH) begin
               // HH high
               digit = (hh/10)%10;
               digit_n = (hh_n/10)%10;
               xofs = (X - FONT_START_X) / FONT_MULTI;
            end else if (FONT_START_X + FONT_WIDTH <= X && X < FONT_START_X + FONT_WIDTH*2) begin
               // HH low
               digit = hh%10;
               digit_n = hh_n%10;
               xofs = (X - (FONT_START_X + FONT_WIDTH)) / FONT_MULTI;
            end else if (FONT_START_X + FONT_WIDTH*2 <= X && X < FONT_START_X + FONT_WIDTH*2 + DOT_WIDTH) begin
               // :
               xofs = (X - (FONT_START_X + FONT_WIDTH*2)) / FONT_MULTI;
`ifdef BLINK_COLON
               if (nframe < 30) begin
                  digit = 10; // colon
                  digit_n = 10;
               end else begin
                  digit = 12; // blank
                  digit_n = 12;
               end
`else
               digit = 10; // colon
               digit_n = 10;
`endif
            end else if (FONT_START_X + FONT_WIDTH*2 + DOT_WIDTH <= X && X < FONT_START_X + FONT_WIDTH*3 + DOT_WIDTH) begin
               // MM high
               digit = (mm/10)%10;
               digit_n = (mm_n/ 10) % 10;
               xofs = (X - (FONT_START_X + FONT_WIDTH*2 + DOT_WIDTH)) / FONT_MULTI;
            end else if (FONT_START_X + FONT_WIDTH*3 + DOT_WIDTH <= X && X < FONT_START_X + FONT_WIDTH*4 + DOT_WIDTH) begin
               // MM low
               digit = mm % 10;
               digit_n = mm_n % 10;
               xofs = (X - (FONT_START_X + FONT_WIDTH*3 + DOT_WIDTH)) / FONT_MULTI;
            end else if (FONT_START_X + FONT_WIDTH*4 + DOT_WIDTH <= X && X < FONT_START_X + FONT_WIDTH*4 + DOT_WIDTH*2) begin
               // :
               xofs = (X - (FONT_START_X + FONT_WIDTH*4 + DOT_WIDTH)) / FONT_MULTI;
`ifdef BLINK_COLON
               if (nframe < 30) begin
                  digit = 10; // colon
                  digit_n = 10;
               end else begin
                  digit = 12; // blank
                  digit_n = 12;
               end
`else
               digit = 10; // colon
               digit_n = 10;
`endif
            end else if (FONT_START_X + FONT_WIDTH*4 + DOT_WIDTH*2<= X && X < FONT_START_X + FONT_WIDTH*5 + DOT_WIDTH*2) begin
               // SS high
               digit = (ss/10)%10;
               digit_n = (ss_n/ 10) % 10;
               xofs = (X - (FONT_START_X + FONT_WIDTH*4 + DOT_WIDTH*2)) / FONT_MULTI;
            end else if (FONT_START_X + FONT_WIDTH*5 + DOT_WIDTH*2<= X && X < FONT_START_X + FONT_WIDTH*6 + DOT_WIDTH*2) begin
               // SS low
               digit = ss % 10;
               digit_n = ss_n % 10;
               xofs = (X - (FONT_START_X + FONT_WIDTH*5 + DOT_WIDTH*2)) / FONT_MULTI;
            end else begin
               digit = 12; // none
               digit_n = 12;
            end
         end else begin
            digit = 12;
            digit_n = 12;
         end //

         if (digit != digit_n && 0 <= digit && digit <= 12) begin
            {s[0],s[1],s[2],s[3]} = font_rle(digit, yofs);
            {s[0],s[1],s[2],s[3]} = rle_to_endpoints(s[0],s[1],s[2],s[3]);
            {f[0],f[1],f[2],f[3]} = font_rle(digit_n, yofs);
            {f[0],f[1],f[2],f[3]} = rle_to_endpoints(f[0],f[1],f[2],f[3]);
            {ep[0],ep[1],ep[2],ep[3]} = blend_endpoints(s[0],s[1],s[2],s[3],f[0],f[1],f[2],f[3],nframe);
         end else begin
            {s[0],s[1],s[2],s[3]} = font_rle(digit, yofs);
            {ep[0],ep[1],ep[2],ep[3]} = rle_to_endpoints(s[0],s[1],s[2],s[3]);
         end
         if (ep[0] && ((ep[0] <= xofs && xofs < ep[1]) || (ep[3] != 0 && ep[2] <= xofs && xofs < ep[3]))) begin
            {r_R,r_B,r_G} <= {8'hff,8'hff,8'hff};
         end else begin
            {r_R,r_B,r_G} <= {8'h00,8'h00,8'h00};
         end
      end else begin // if (den)
         {r_R,r_B,r_G} <= {8'h00,8'h00,8'h00};
      end // else: !if(den)

   end // always@ (posedge clk_lcd)

   //
   
   assign R = r_R;
   assign G = r_G;
   assign B = r_B;

endmodule
